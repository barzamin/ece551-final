`default_nettype none
/*------------------------------------------------------------------------------
--  This testbench measures the time it takes for pitch/roll/yaw to converge
--  to a new value at one thrust level, then checks that at 
--  a higher thrust levels the time to converge is smaller.
--
--  Team: MEI
--  Authors:
--    * Mitchell Kitzinger
--    * Erin Marshall
--    * Isaac Colbert
--  Term: Spring 2021
------------------------------------------------------------------------------*/
module QuadCopter_varied_thrust_tb();

endmodule